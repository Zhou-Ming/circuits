.model emitter_tline ltra r=40.35 g=0 l=3.874e-07 c=8.858e-11 len=2.5e-04
