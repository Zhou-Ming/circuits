.model emitter_tline ltra r=42.2 g=0 l=2.567e-07 c=1.442e-10 len=4.45e-04
